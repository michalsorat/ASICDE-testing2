module rootModule500_sa0_0_sa1_0();
    rootModule500_sa0_0_sa1_0_sa2_0 inst_0();
endmodule
