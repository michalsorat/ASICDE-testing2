module rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0();
    rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0 inst_0();
endmodule
