module rootModule400_sa0_0();
    rootModule400_sa0_0_sa1_0 inst_0();
endmodule
