module rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0();
    rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0 inst_0();
    rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_1 inst_1();
    rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_2 inst_2();
    rootModule500_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_3 inst_3();
endmodule
