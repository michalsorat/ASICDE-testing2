module rootModule1000_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0();
    rootModule1000_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0 inst_0();
endmodule
