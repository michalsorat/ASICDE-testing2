module rootModule1000_sa0_0_sa1_0_sa2_0_sa3_0();
    rootModule1000_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0 inst_0();
endmodule
