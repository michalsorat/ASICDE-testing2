module rootModule400_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_2_sa7_0_sa8_2_sa9_1();
endmodule
