module rootModule1000_sb0_0_sb1_0_sb2_0();
    rootModule1000_sb0_0_sb1_0_sb2_0_sb3_0 inst_0();
endmodule
