module rootModule1000_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_1_sb8_3_sb9_4();
endmodule
