module rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_4_sa8_0_sa9_3();
endmodule
