module rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1();
    rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1_sa9_0 inst_0();
    rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1_sa9_1 inst_1();
    rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1_sa9_2 inst_2();
    rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1_sa9_3 inst_3();
    rootModule200_sa0_0_sa1_0_sa2_0_sa3_0_sa4_0_sa5_0_sa6_0_sa7_3_sa8_1_sa9_4 inst_4();
endmodule
