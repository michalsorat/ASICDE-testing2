module rootModule200_sa0_0();
    rootModule200_sa0_0_sa1_0 inst_0();
endmodule
