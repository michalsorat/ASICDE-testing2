module rootModule1000();
    rootModule1000_sa0_0 inst_0();
endmodule
