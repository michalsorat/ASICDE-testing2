module rootModule1000_sa0_0_sa1_0();
    rootModule1000_sa0_0_sa1_0_sa2_0 inst_0();
endmodule
