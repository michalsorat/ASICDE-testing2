module rootModule500();
    rootModule500_sa0_0 inst_0();
endmodule
