module rootModule200();
    rootModule200_sa0_0 inst_0();
endmodule
