module rootModule400();
    rootModule400_sa0_0 inst_0();
endmodule
