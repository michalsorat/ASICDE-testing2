module rootModule1000();
    rootModule1000_sb0_0 inst_0();
endmodule
