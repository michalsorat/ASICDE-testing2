module rootModule1000_sb0_0();
    rootModule1000_sb0_0_sb1_0 inst_0();
endmodule
